--------------------------------------------------------------------------------
-- Synthesizer : ISE 14.6
-- Platform    : Linux Ubuntu 10.04
-- Targets     : Synthese
--------------------------------------------------------------------------------
-- This work is held in copyright as an unpublished work by HEPHY (Institute
-- of High Energy Physics) All rights reserved.  This work may not be used
-- except by authorized licensees of HEPHY. This work is the
-- confidential information of HEPHY.
--------------------------------------------------------------------------------
-- $HeadURL: svn://heros.hephy.oeaw.ac.at/GlobalTriggerUpgrade/firmware/uGT_fw_integration/trunk/uGT_algos/firmware/hdl/gt_mp7_top_pkg_tpl.vhd $
-- $Date: 2015-05-21 15:33:04 +0200 (Thu, 21 May 2015) $
-- $Author: wittmann $
-- $Revision: 3966 $
--------------------------------------------------------------------------------
--
-- Notes on using `gtu-pkgpatch-ipbus' for this package:
--  * {{IPBUS_TIMESTAMP}}    32 bit UNIX timestamp placeholder (X"00000000")
--  * {{IPBUS_USERNAME}}     unix username 32 char string placeholder (X"...")
--  * {{IPBUS_HOSTNAME}}     machine hostname 32 char string placeholder (X"...")
--  * {{IPBUS_BUILD_VERSION}}     build firmware version (X"...")
--
--------------------------------------------------------------------------------

-- HB 2016-06-30: removed unused constants and comments

library IEEE;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use work.mp7_brd_decl.all;

package gt_mp7_top_pkg is

-- BA 2014-08-06: TIMESTAMP generated by gtu-pkgpatch-ipbus (32 bits), has to be interpreted as 32 bit UNIX timestamp.
constant TOP_TIMESTAMP : std_logic_vector(31 downto 0) := X"5b8f8fb9";
-- HB 2014-05-23: USERNAME generated by gtu-pkgpatch-ipbus (256 bits = 8 x 32 bits), has to be interpreted as 32 ASCII-characters string (from right to left).
constant TOP_USERNAME : std_logic_vector(32*8-1 downto 0)  := X"0000000000000000000000000000000000000000000000007265756167726562";
-- HB 2014-05-23: HOSTNAME generated by gtu-pkgpatch-ipbus (256 bits = 8 x 32 bits), has to be interpreted as 32 ASCII-characters string (from right to left).
constant TOP_HOSTNAME : std_logic_vector(32*8-1 downto 0) := X"000000000000000000000000000000000000000000000068746e79732d746775";
-- JW 2015-05-21: TOP_VERSION generated by gtu-pkgpatch-ipbus (32 bits), is the overall version number for a gt_mp7 build (e.g. 1003 for v1003)
constant TOP_BUILD_VERSION : std_logic_vector(31 downto 0) := X"00008106";

end;



